/*************************************************
*
* This CDL file subfsa_eod.cdl was created with cfgedit
* version 6.0.01
*
**************************************************/

bindArch AuRA.naval;

[
FSA1:FSA(
      society[$AN_2821]<809,279>|State2| = [
          %Objects = {Mines},
          %move_to_object_gain = {1.0},
          %avoid_obstacle_gain = {1.0},
          %wander_gain = {0.0},
          %avoid_obstacle_sphere = {2.2},
          %avoid_obstacle_safety_margin = {0.3}
,
        MoveToward]<100,100>
,
      society[$AN_2823]<810,492>|State3| = [
        Stop]<100,100>
,
      society[$AN_2825]<541,493>|State5| = [
          %Object = {Mine}
,
        TerminateObject]<100,100>
,
      society[$AN_2827]<256,491>|State6| = [
          %notify_message = {"EODTask completed."}
,
        Notify]<100,100>
,
      society[Start]<50,50>|Start| = [
        Stop]<100,100>
,
      society[$AN_2830]<258,669>|State7| = [
        Stop]<10,10>
,
      society[$AN_2832]<424,115>|State8| = [
          %move_to_object_gain = {1.0},
          %avoid_obstacle_gain = {1.0},
          %wander_gain = {0.0},
          %avoid_obstacle_sphere = {2.2},
          %avoid_obstacle_safety_margin = {0.3}
,
        MoveToward_NotifiedObject]<10,10>
,
      society[$AN_2834]<595,279>|State9| = [
        Stop]<10,10>
,
      society[$AN_2836]<256,278>|State1| = [
        Stop]<100,100>
,
      society[$AN_2858]<808,108>|State9| = [
          %Objects = {Friendly_Robots},
          %move_away_object_gain = {1.0},
          %avoid_obstacle_gain = {0.5},
          %wander_gain = {0.0},
          %avoid_objects_sphere = {100.0},
          %avoid_objects_safety_margin = {10.0},
          %avoid_obstacle_sphere = {1.2},
          %avoid_obstacle_safety_margin = {0.3}
,
        MoveAway]<10,10>
,
      rules[$AN_2836]<256,278>|State1| = if [
          %Objects = {Mines}
,
        NotDetected]<0,0>|Trans8|
 goto $AN_2827,
      rules[Start]<50,50>|Start| = if [
        Immediate]<0,0>|Trans1|
 goto $AN_2836,
      rules[$AN_2827]<256,491>|State6| = if [
        Immediate]<0,0>|Trans1|
 goto $AN_2830,
      rules[$AN_2825]<541,493>|State5| = if [
          %Delay = {1.0}
,
        Wait]<411,493>|Trans7|
 goto $AN_2827,
      rules[$AN_2834]<595,279>|State9| = if [
          %Objects = {Mines}
,
        Detect]<0,0>|Trans2|
 goto $AN_2821,
      rules[$AN_2836]<256,278>|State1| = if [
          %Delay = {5.0}
,
        Wait]<0,0>|Trans2|
 goto $AN_2834,
      rules[$AN_2836]<256,278>|State1| = if [
        Notified_ObjectLocation]<0,0>|Trans3|
 goto $AN_2832,
      rules[$AN_2821]<809,279>|State2| = if [
          %Objects = {Mines},
          %Distance = {20.0}
,
        Near]<0,0>|Trans3|
 goto $AN_2823,
      rules[$AN_2823]<810,492>|State3| = if [
          %Delay = {1.0}
,
        Wait]<0,0>|Trans6|
 goto $AN_2825,
      rules[$AN_2832]<424,115>|State8| = if [
          %Distance = {20}
,
        NearNotifiedObject]<0,0>|Trans6|
 goto $AN_2834,
      rules[$AN_2821]<809,279>|State2| = if [
          %Objects = {Friendly_Robots},
          %Distance = {50.0}
,
        Near]<0,0>|Trans1|
 goto $AN_2858,
      rules[$AN_2858]<808,108>|State9| = if [
          %Objects = {Friendly_Robots},
          %Distance = {60.0}
,
        AwayFrom]<0,0>|Trans2|
 goto $AN_2821)<33,49>|The State Machine|
]<10,10>

