/*************************************************
*
* This CDL file preserve.cdl was created with cfgedit
* version 6.0.01
*
**************************************************/

bindArch AuRA.urban;

instBP<227,266> $AN_1579 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1588,
            rules[$AN_1588]<199,330>|State1| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1591,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1588]<199,330>|State1| = [
              InitiaizeCSB]<100,100>
,
            society[$AN_1591]<588,328>|State2| = [
              UpdateCSBSensorData]<100,100>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1595 from movement(
  base_vel = {0.1},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[$AN_1610]<594,264>|State3| = [
              Stop]<100,100>
,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1613]<241,268>|State1| = [
              Standby*]<100,100>
,
            society[$AN_1615]<724,606>|State2| = [
                %method = {Comm_Preserve},
                %follow_csb_advise_gain = {1.0},
                %avoid_obstacle_gain = {0.04},
                %wander_gain = {0.0},
                %avoid_obstacle_sphere = {4.0},
                %avoid_obstacle_safety_margin = {0.5}
,
              FollowCSBAdvise]<100,100>
,
            society[$AN_1617]<241,602>|State4| = [
                %Goal_Location = {119.0, 33.0},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.03},
                %avoid_obstacle_sphere = {1.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1749]<727,895>|State5| = [
              Stop]<10,10>
,
            rules[$AN_1613]<241,268>|State1| = if [
                %notify_message = {"MOTOR FAILURE DETECTED"}
,
              TaskExited]<0,0>|Trans2|
 goto $AN_1610,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans19|
 goto $AN_1613,
            rules[$AN_1613]<241,268>|State1| = if [
                %notify_message = {"PROCEED MISSION"}
,
              TaskExited]<0,0>|Trans1|
 goto $AN_1617,
            rules[$AN_1617]<241,602>|State4| = if [
                %Goal_Tolerance = {0.5},
                %Goal_Location = {119.0, 33.0}
,
              AtGoal]<0,0>|Trans2|
 goto $AN_1615,
            rules[$AN_1615]<724,606>|State2| = if [
                %notify_message = {"Mission Accomplished"}
,
              Notified]<0,0>|Trans6|
 goto $AN_1749)<292,156>|The State Machine|
,
        max_vel = {1.6},
        base_vel = {1.4},
        cautious_vel = {0.3},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<100,100> $AN_1627 from vehicle(
  bound_to = preserveRobot3:DEFAULT_ROBOT(
preserveRobot3:[
          $AN_1595,
          $AN_1579]
)<22,348>|Individual Robot|
);

instBP<227,266> $AN_1628 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1588,
            rules[$AN_1588]<199,330>|State1| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1591,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1588]<199,330>|State1| = [
              InitiaizeCSB]<100,100>
,
            society[$AN_1591]<588,328>|State2| = [
              UpdateCSBSensorData]<100,100>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1642 from movement(
  base_vel = {0.1},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[$AN_1610]<594,264>|State3| = [
              Stop]<100,100>
,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1613]<241,268>|State1| = [
              Standby*]<100,100>
,
            society[$AN_1660]<1020,600>|State4| = [
                %Goal_Location = {126.5, 32.5},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.03},
                %avoid_obstacle_sphere = {1.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1662]<570,600>|State5| = [
                %Goal_Location = {147.5, 48.0},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.03},
                %avoid_obstacle_sphere = {1.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1664]<115,600>|State6| = [
                %Goal_Location = {130.0, 51.0},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.03},
                %avoid_obstacle_sphere = {1.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1666]<1021,986>|State6| = [
                %Goal_Location = {135.0, 72.0},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.03},
                %avoid_obstacle_sphere = {1.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1668]<597,982>|State7| = [
                %Goal_Location = {141.0, 98.0},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.03},
                %avoid_obstacle_sphere = {1.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1670]<132,982>|State8| = [
                %Goal_Location = {141.0, 104.0},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.03},
                %avoid_obstacle_sphere = {1.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1672]<131,1345>|State9| = [
                %Goal_Location = {141.0, 98.0},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.03},
                %avoid_obstacle_sphere = {1.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1729]<630,1354>|State10| = [
                %Goal_Location = {135.0, 72.0},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.03},
                %avoid_obstacle_sphere = {1.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1733]<1017,1359>|State11| = [
                %Goal_Location = {130.0, 51.0},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.03},
                %avoid_obstacle_sphere = {1.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1737]<1021,1675>|State12| = [
              Stop]<10,10>
,
            society[$AN_1741]<616,1674>|State13| = [
                %notify_message = {"Mission Accomplished"}
,
              NotifyRobots]<10,10>
,
            society[$AN_1745]<213,1677>|State14| = [
              Stop]<10,10>
,
            rules[$AN_1613]<241,268>|State1| = if [
                %notify_message = {"MOTOR FAILURE DETECTED"}
,
              TaskExited]<0,0>|Trans2|
 goto $AN_1610,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans19|
 goto $AN_1613,
            rules[$AN_1660]<1020,600>|State4| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {126.5, 32.5}
,
              AtGoal]<812,657>|Trans1|
 goto $AN_1662,
            rules[$AN_1662]<570,600>|State5| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {147.5, 48.0}
,
              AtGoal]<0,0>|Trans2|
 goto $AN_1664,
            rules[$AN_1666]<1021,986>|State6| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {135.0, 72.0}
,
              AtGoal]<0,0>|Trans5|
 goto $AN_1668,
            rules[$AN_1668]<597,982>|State7| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {141.0, 98.0}
,
              AtGoal]<0,0>|Trans6|
 goto $AN_1670,
            rules[$AN_1670]<132,982>|State8| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {141.0, 104.0}
,
              AtGoal]<0,0>|Trans7|
 goto $AN_1672,
            rules[$AN_1613]<241,268>|State1| = if [
                %notify_message = {"PROCEED MISSION"}
,
              TaskExited]<585,414>|Trans1|
 goto $AN_1660,
            rules[$AN_1664]<115,600>|State6| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {130.0, 51.0}
,
              AtGoal]<10,10>|Trans9|
 goto $AN_1666,
            rules[$AN_1672]<131,1345>|State9| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {141.0, 98.0}
,
              AtGoal]<0,0>|Trans1|
 goto $AN_1729,
            rules[$AN_1729]<630,1354>|State10| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {135.0, 72.0}
,
              AtGoal]<10,10>|Trans2|
 goto $AN_1733,
            rules[$AN_1733]<1017,1359>|State11| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {130.0, 51.0}
,
              AtGoal]<0,0>|Trans3|
 goto $AN_1737,
            rules[$AN_1737]<1021,1675>|State12| = if [
                %Delay = {10.0}
,
              Wait]<0,0>|Trans4|
 goto $AN_1741,
            rules[$AN_1741]<616,1674>|State13| = if [
              MessageSent]<0,0>|Trans5|
 goto $AN_1745)<292,156>|The State Machine|
,
        max_vel = {1.6},
        base_vel = {1.4},
        cautious_vel = {0.3},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<100,100> $AN_1692 from vehicle(
  bound_to = preserveRobot2:DEFAULT_ROBOT(
preserveRobot2:[
          $AN_1642,
          $AN_1628]
)<22,190>|Individual Robot|
);

instBP<227,266> $AN_1693 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1588,
            rules[$AN_1588]<199,330>|State1| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1591,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1588]<199,330>|State1| = [
              InitiaizeCSB]<100,100>
,
            society[$AN_1591]<588,328>|State2| = [
              UpdateCSBSensorData]<100,100>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1707 from movement(
  base_vel = {0.1},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1610]<229,284>|State3| = [
              Stop]<100,100>
,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans2|
 goto $AN_1610)<292,156>|The State Machine|
,
        max_vel = {1.6},
        base_vel = {1.4},
        cautious_vel = {0.3},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<120,120> $AN_1726 from vehicle(
  bound_to = preserveRobot1:DEFAULT_ROBOT(
preserveRobot1:[
          $AN_1707,
          $AN_1693]
)<22,36>|Individual Robot|
);

[
[
    $AN_1726,
    $AN_1692,
    $AN_1627]<10,10>|Group of Robots|
]<10,10>

