/*************************************************
*
* This CDL file sample_inspect.cdl was created with cfgedit
* version 6.0.01
*
**************************************************/

bindArch AuRA.naval;

instBP<222,15> |The Wheels Binding Point| $AN_2376 from movement(
  base_vel = {2.5},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA1:FSA(
            society[Start]<50,50>|Start| = [
              Stop]<10,10>
,
            society[$AN_2391]<299,273>|State1| = [
              Stop]<10,10>
,
            society[$AN_2393]<662,275>|State2| = [
                %Objects = {Enemies},
                %move_to_object_gain = {1.0},
                %avoid_obstacle_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_sphere = {2.2},
                %avoid_obstacle_safety_margin = {0.3}
,
              MoveToward]<10,10>
,
            society[$AN_2395]<661,503>|State3| = [
                %notify_message = {"Enemy put down weapons."}
,
              NotifyRobots]<10,10>
,
            society[$AN_2397]<312,501>|State4| = [
              Stop]<10,10>
,
            society[$AN_2399]<311,712>|State5| = [
                %Objects = {Illegal_Weapons}
,
              LookFor]<10,10>
,
            society[$AN_2401]<309,975>|State6| = [
                %alert_subject = {"Warning: Illegal weapons seized"},
                %alert_message = {"The robot has found illegal weapons."},
                %sends_email = {NO_Email},
                %recipient = {""},
                %sends_image = {NO_Image}
,
              Alert]<10,10>
,
            society[$AN_2403]<693,852>|State7| = [
                %alert_subject = {"Warning: No weapon found"},
                %alert_message = {""},
                %sends_email = {NO_Email},
                %recipient = {""},
                %sends_image = {NO_Image}
,
              Alert]<10,10>
,
            society[$AN_2405]<696,1069>|State8| = [
              Stop]<10,10>
,
            rules[$AN_2391]<299,273>|State1| = if [
                %notify_message = {"Enemy stop."}
,
              Notified]<477,275>|Trans2|
 goto $AN_2393,
            rules[$AN_2393]<662,275>|State2| = if [
                %Objects = {Enemies},
                %Distance = {5.0}
,
              Near]<0,0>|Trans3|
 goto $AN_2395,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_2391,
            rules[$AN_2395]<661,503>|State3| = if [
              MessageSent]<10,10>|Trans5|
 goto $AN_2397,
            rules[$AN_2397]<312,501>|State4| = if [
                %Delay = {1.0}
,
              Wait]<0,0>|Trans6|
 goto $AN_2399,
            rules[$AN_2399]<311,712>|State5| = if [
                %Objects = {Illegal_Weapons},
                %Distance = {30.0}
,
              Near]<312,804>|Trans7|
 goto $AN_2401,
            rules[$AN_2399]<311,712>|State5| = if [
                %Delay = {3.0}
,
              Wait]<516,788>|Trans8|
 goto $AN_2403,
            rules[$AN_2401]<309,975>|State6| = if [
              Alerted]<10,10>|Trans9|
 goto $AN_2405,
            rules[$AN_2403]<693,852>|State7| = if [
              Alerted]<10,10>|Trans10|
 goto $AN_2405)<292,156>|The State Machine|
,
        max_vel = {5.0},
        base_vel = {2.5},
        cautious_vel = {0.5},
        cautious_mode = {false})<222,15>|The Wheel Actuator|
);

instBP<0,0> $AN_2425 from vehicle(
  bound_to = sample_inspectRobot1:DEFAULT_ROBOT(
sample_inspectRobot1:[
          $AN_2376]
)<0,0>|Individual Robot|
);

[
[
    $AN_2425]<10,10>|Group of Robots|
]<10,10>

