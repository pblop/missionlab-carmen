/*************************************************
*
* This CDL file /hr7/projects/robot/mission/src/usability_demos/Task0/example.cdl was created with cfgedit
* version 1.0a
*
**************************************************/

bindArch AuRA;

instGroup $AN_221 from [
    %Objects = {Mines}
,
  PickUp];
instGroup $AN_222 from [
    %Objects = {Mines}
,
  MoveTo];
instGroup $AN_223 from [
  Stop];
instBP<565,111> |The Wheels Binding Point| $AN_224 from movement(
  v<0,0> = ,
  base_vel = {0.1},
  bound_to = base:DRIVE(
        v<292,156> = FSA(
            society[Start]<135,192>|Start| = $AN_223,
            society[$AN_240]<372,195>|State1| = $AN_222,
            society[$AN_244]<692,222>|State2| = $AN_221,
            society[$AN_252]<374,438>|State3| = [
              Stop]<10,10>
,
            rules[$AN_240]<372,195>|State1| = if [
                %Objects = {Mines},
                %Distance = {0.2}
,
              Near]<546,252>|Trans2|
 goto $AN_244,
            rules[$AN_244]<692,222>|State2| = if [
              FirstTime]<10,10>|Trans3|
 goto $AN_240,
            rules[Start]<135,192>|Start| = if [
              FirstTime]<0,0>|Trans1|
 goto $AN_240,
            rules[$AN_240]<372,195>|State1| = if [
                %Objects = {Mines}
,
              UnDetect]<0,0>|Trans1|
 goto $AN_252)<292,156>|The State Machine|
,
        max_vel = {0.2},
        base_vel = {1},
        cautious_vel = {0.05},
        cautious_mode = {false})<565,111>|The Wheels Actuator|
);

instBP<0,0> $AN_303 from vehicle(
  bound_to = exampleRobot1:MRV2(
exampleRobot1:[
          $AN_224]
)<0,0>|The robot|
);

[
[
    $AN_303]<0,0>|The Configuration|
]<10,10>
