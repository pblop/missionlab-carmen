/*************************************************
*
* This CDL file testCMDLi-single.cdl was created with cfgedit
* version 6.0.01
*
**************************************************/

bindArch AuRA.urban;

instBP<227,266> $AN_1620 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<10,10>|Trans1|
 goto $AN_1590,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1590]<195,164>|State1| = [
              Stop]<10,10>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1631 from movement(
  v<0,0> = ,
  base_vel = {0.1},
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[Start]<50,50>|Start| = [
              Stop]<10,10>
,
            society[$AN_1610]<208,211>|State2| = [
              Standby*]<10,10>
,
            society[$AN_1611]<572,215>|State3| = [
                %env_filename = {"TSRB_Parking-8F.ovl"},
                %cmdl_filename = {"testCMDLi-single.cmdl"},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.0},
                %avoid_obstacle_sphere = {3.0},
                %avoid_obstacle_safety_margin = {0.5},
                %goal_tolerance = {1.0}
,
              FollowCMDLiCommands]<10,10>
,
            society[$AN_1612]<210,455>|State4| = [
              Stop]<10,10>
,
            rules[$AN_1610]<208,211>|State2| = if [
                %notify_message = {"PROCEED MISSION"}
,
              TaskExited]<0,0>|Trans1|
 goto $AN_1611,
            rules[$AN_1610]<208,211>|State2| = if [
                %notify_message = {"MOTOR FAILURE DETECTED"}
,
              TaskExited]<0,0>|Trans2|
 goto $AN_1612,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans3|
 goto $AN_1610)<292,156>|The State Machine|
,
        max_vel = {1.6},
        base_vel = {1.4},
        cautious_vel = {0.7},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<0,0> $AN_1656 from vehicle(
  bound_to = testCMDLi-singleRobot1:DEFAULT_ROBOT(
testCMDLi-singleRobot1:[
          $AN_1631,
          $AN_1620]
)<35,29>|Individual Robot|
);

[
[
    $AN_1656]<10,10>|Group of Robots|
]<10,10>

