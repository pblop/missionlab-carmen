/*************************************************
*
* This CDL file sample_cbr_behavioral_select.cdl was created with cfgedit
* version 5.0.08
*
**************************************************/

bindArch AuRA.urban;

instBP<227,266> $AN_1508 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<10,10>|Trans1|
 goto $AN_1517,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1517]<195,164>|State1| = [
              Stop]<10,10>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1520 from movement(
  base_vel = {0.1},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[Start]<50,50>|Start| = [
              Stop]<10,10>
,
            society[$AN_1536]<321,250>|State1| = [
                %Goal_Location = {71, 30},
                %avoid_obstacle_gain = {0.5},
                %obstacle_safety_margin = {0.75}
,
              GoToOutdoor_CBR]<10,10>
,
            society[$AN_1538]<759,117>|State2| = [
                %load_new_overlay = {DEFAULT_MAP},
                %new_overlay = {"Empty.ovl"}
,
              ResetWorld]<10,10>
,
            rules[Start]<50,50>|Start| = if [
              Immediate]<10,10>|Trans1|
 goto $AN_1536,
            rules[$AN_1536]<321,250>|State1| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {71, 30}
,
              AtGoal]<10,10>|Trans1|
 goto $AN_1538)<292,156>|The State Machine|
,
        max_vel = {0.6},
        base_vel = {0.5},
        cautious_vel = {0.3},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<0,0> $AN_1544 from vehicle(
  bound_to = sample_cbr_behavioral_selectRobot1:DEFAULT_ROBOT(
sample_cbr_behavioral_selectRobot1:[
          $AN_1520,
          $AN_1508]
)<0,0>|Individual Robot|
);

NoName:[
[
    $AN_1544]<10,10>|Group of Robots|
]<10,10>

