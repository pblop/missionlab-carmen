/*************************************************
*
* This CDL file tsrb-bnf.cdl was created with cfgedit
* version 6.0.01
*
**************************************************/

bindArch AuRA.urban;

instBP<227,266> $AN_1596 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<10,10>|Trans1|
 goto $AN_1605,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1605]<195,164>|State1| = [
              Stop]<10,10>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1608 from movement(
  v<0,0> = ,
  base_vel = {0.1},
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[Start]<50,50>|Start| = [
              Stop]<10,10>
,
            society[$AN_1627]<120,300>|State1| = [
                %Goal_Location = {13.18, 13.50},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.0},
                %avoid_obstacle_sphere = {2.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1629]<752,312>|State2| = [
                %Goal_Location = {14.11, 29.89},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.0},
                %avoid_obstacle_sphere = {2.5},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            rules[$AN_1627]<120,300>|State1| = if [
                %Goal_Tolerance = {2.0},
                %Goal_Location = {13.18, 13.50}
,
              AtGoal]<0,0>|Trans4|
 goto $AN_1629,
            rules[Start]<50,50>|Start| = if [
              Immediate]<10,10>|Trans5|
 goto $AN_1627,
            rules[$AN_1629]<752,312>|State2| = if [
                %Goal_Tolerance = {2.0},
                %Goal_Location = {14.11, 29.89}
,
              AtGoal]<0,0>|Trans6|
 goto $AN_1627)<292,156>|The State Machine|
,
        max_vel = {2.0},
        base_vel = {1.5},
        cautious_vel = {0.05},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<0,0> $AN_1624 from vehicle(
  bound_to = tsrb-bnfRobot1:DEFAULT_ROBOT(
tsrb-bnfRobot1:[
          $AN_1608,
          $AN_1596]
)<0,0>|Individual Robot|
);

[
[
    $AN_1624]<10,10>|Group of Robots|
]<10,10>

