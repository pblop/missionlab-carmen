/*************************************************
*
* This CDL file sample_CSB2.cdl was created with cfgedit
* version 6.0.01
*
**************************************************/

bindArch AuRA.urban;

instBP<227,266> $AN_1555 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1564,
            rules[$AN_1564]<199,330>|State1| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1567,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1564]<199,330>|State1| = [
              InitiaizeCSB]<100,100>
,
            society[$AN_1567]<588,328>|State2| = [
              UpdateCSBSensorData]<100,100>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1571 from movement(
  base_vel = {0.1},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1587]<220,381>|State1| = [
                %method = {Internalized_Plan},
                %follow_csb_advise_gain = {1.0},
                %avoid_obstacle_gain = {0.5},
                %wander_gain = {0.0},
                %avoid_obstacle_sphere = {1.2},
                %avoid_obstacle_safety_margin = {0.3}
,
              FollowCSBAdvise]<100,100>
,
            society[$AN_1589]<753,396>|State3| = [
                %method = {Comm_Recovery},
                %follow_csb_advise_gain = {1.0},
                %avoid_obstacle_gain = {0.5},
                %wander_gain = {0.0},
                %avoid_obstacle_sphere = {1.2},
                %avoid_obstacle_safety_margin = {0.3}
,
              FollowCSBAdvise]<100,100>
,
            society[$AN_1635]<499,194>|State3| = [
                %alert_subject = {"Weak Signal!"},
                %alert_message = {"The robot is now trying to recover communication."},
                %sends_email = {NO_Email},
                %recipient = {""},
                %sends_image = {NO_Image}
,
              Alert]<10,10>
,
            society[$AN_1643]<496,544>|State4| = [
                %alert_subject = {"Communication Recovered!"},
                %alert_message = {"The robot is now resuming the internalized plan."},
                %sends_email = {NO_Email},
                %recipient = {""},
                %sends_image = {NO_Image}
,
              Alert]<10,10>
,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans2|
 goto $AN_1587,
            rules[$AN_1587]<220,381>|State1| = if [
                %threshold = {35.0}
,
              WeakCommSignal]<0,0>|Trans2|
 goto $AN_1635,
            rules[$AN_1635]<499,194>|State3| = if [
              Alerted]<0,0>|Trans2|
 goto $AN_1589,
            rules[$AN_1589]<753,396>|State3| = if [
                %threshold = {45.0}
,
              StrongCommSignal]<650,457>|Trans1|
 goto $AN_1643,
            rules[$AN_1643]<496,544>|State4| = if [
              Alerted]<10,10>|Trans4|
 goto $AN_1587)<292,156>|The State Machine|
,
        max_vel = {1.6},
        base_vel = {1.4},
        cautious_vel = {0.7},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<100,100> $AN_1597 from vehicle(
  bound_to = sample_CSB2Robot2:DEFAULT_ROBOT(
sample_CSB2Robot2:[
          $AN_1571,
          $AN_1555]
)<28,200>|Individual Robot|
);

instBP<227,266> $AN_1598 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1564,
            rules[$AN_1564]<199,330>|State1| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1567,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1564]<199,330>|State1| = [
              InitiaizeCSB]<10,10>
,
            society[$AN_1567]<588,328>|State2| = [
              UpdateCSBSensorData]<10,10>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1612 from movement(
  base_vel = {0.1},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[Start]<50,50>|Start| = [
              Stop]<10,10>
,
            society[$AN_1628]<240,267>|State1| = [
                %method = {Internalized_Plan},
                %follow_csb_advise_gain = {1.0},
                %avoid_obstacle_gain = {0.5},
                %wander_gain = {0.0},
                %avoid_obstacle_sphere = {1.2},
                %avoid_obstacle_safety_margin = {0.3}
,
              FollowCSBAdvise]<10,10>
,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans19|
 goto $AN_1628)<292,156>|The State Machine|
,
        max_vel = {1.6},
        base_vel = {1.4},
        cautious_vel = {0.7},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<0,0> $AN_1632 from vehicle(
  bound_to = sample_CSB2Robot1:DEFAULT_ROBOT(
sample_CSB2Robot1:[
          $AN_1612,
          $AN_1598]
)<27,38>|Individual Robot|
);

[
[
    $AN_1632,
    $AN_1597]<10,10>|Group of Robots|
]<10,10>

