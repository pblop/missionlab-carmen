/*************************************************
*
* This CDL file tsrb-bnf2-oa-off.cdl was created with cfgedit
* version 6.0.01
*
**************************************************/

bindArch AuRA.urban;

instBP<227,266> $AN_1555 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<10,10>|Trans1|
 goto $AN_1564,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1564]<195,164>|State1| = [
              Stop]<10,10>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1567 from movement(
  v<0,0> = ,
  base_vel = {0.1},
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[Start]<50,50>|Start| = [
              Stop]<10,10>
,
            society[$AN_1583]<734,368>|State1| = [
                %Goal_Location = {53.08, 37.432},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.0},
                %avoid_obstacle_sphere = {5.0},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            society[$AN_1585]<156,362>|State2| = [
                %Goal_Location = {62.08, 37.432},
                %move_to_location_gain = {1.0},
                %wander_gain = {0.0},
                %avoid_obstacle_gain = {0.0},
                %avoid_obstacle_sphere = {5.0},
                %avoid_obstacle_safety_margin = {0.5}
,
              GoTo]<10,10>
,
            rules[Start]<50,50>|Start| = if [
              Immediate]<10,10>|Trans2|
 goto $AN_1585,
            rules[$AN_1585]<156,362>|State2| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {62.08, 37.432}
,
              AtGoal]<0,0>|Trans3|
 goto $AN_1583,
            rules[$AN_1583]<734,368>|State1| = if [
                %Goal_Tolerance = {1.0},
                %Goal_Location = {53.08, 37.432}
,
              AtGoal]<0,0>|Trans4|
 goto $AN_1585)<292,156>|The State Machine|
,
        max_vel = {2.0},
        base_vel = {1.75},
        cautious_vel = {0.05},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<0,0> $AN_1593 from vehicle(
  bound_to = tsrb-bnf2-oa-offRobot1:DEFAULT_ROBOT(
tsrb-bnf2-oa-offRobot1:[
          $AN_1567,
          $AN_1555]
)<0,0>|Individual Robot|
);

[
[
    $AN_1593]<10,10>|Group of Robots|
]<10,10>

