/*************************************************
*
* This CDL file sample_CSB.cdl was created with cfgedit
* version 6.0.01
*
**************************************************/

bindArch AuRA.urban;

instBP<227,266> $AN_1555 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1564,
            rules[$AN_1564]<199,330>|State1| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1567,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1564]<199,330>|State1| = [
              InitiaizeCSB]<100,100>
,
            society[$AN_1567]<588,328>|State2| = [
              UpdateCSBSensorData]<100,100>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1571 from movement(
  v<0,0> = ,
  base_vel = {0.1},
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[$AN_1587]<239,320>|State1| = [
                %method = {Comm_Preserve},
                %follow_csb_advise_gain = {1.0},
                %avoid_obstacle_gain = {0.5},
                %wander_gain = {0.0},
                %avoid_obstacle_sphere = {1.2},
                %avoid_obstacle_safety_margin = {0.3}
,
              FollowCSBAdvise]<100,100>
,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans2|
 goto $AN_1587)<292,156>|The State Machine|
,
        max_vel = {1.6},
        base_vel = {1.4},
        cautious_vel = {0.7},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<100,100> $AN_1605 from vehicle(
  bound_to = sample_CSB2Robot2:DEFAULT_ROBOT(
sample_CSB2Robot2:[
          $AN_1571,
          $AN_1555]
)<28,200>|Individual Robot|
);

instBP<227,266> $AN_1606 from pantilt(
  look_loc<0,0> = ,
  bound_to = camera:PANTILT(
        look_loc<14,299> = FSA(
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1564,
            rules[$AN_1564]<199,330>|State1| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_1567,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_1564]<199,330>|State1| = [
              InitiaizeCSB]<10,10>
,
            society[$AN_1567]<588,328>|State2| = [
              UpdateCSBSensorData]<10,10>
)<11,182>|The State Machine|
)<224,298>|The Camera Actuator|
);

instBP<222,15> |The Wheels Binding Point| $AN_1620 from movement(
  v<0,0> = ,
  base_vel = {0.1},
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA(
            society[Start]<50,50>|Start| = [
              Stop]<10,10>
,
            society[$AN_1636]<240,267>|State1| = [
                %method = {Internalized_Plan},
                %follow_csb_advise_gain = {1.0},
                %avoid_obstacle_gain = {0.5},
                %wander_gain = {0.0},
                %avoid_obstacle_sphere = {1.2},
                %avoid_obstacle_safety_margin = {0.3}
,
              FollowCSBAdvise]<10,10>
,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans19|
 goto $AN_1636)<292,156>|The State Machine|
,
        max_vel = {1.6},
        base_vel = {1.4},
        cautious_vel = {0.7},
        cautious_mode = {true})<222,15>|The Wheel Actuator|
);

instBP<0,0> $AN_1640 from vehicle(
  bound_to = sample_CSB2Robot1:DEFAULT_ROBOT(
sample_CSB2Robot1:[
          $AN_1620,
          $AN_1606]
)<27,38>|Individual Robot|
);

[
[
    $AN_1640,
    $AN_1605]<10,10>|Group of Robots|
]<10,10>

