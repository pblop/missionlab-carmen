/*************************************************
*
* This CDL file sample-type-I-intercept.cdl was created with cfgedit
* version 6.0.01
*
**************************************************/

bindArch AuRA.naval;

instBP<222,15> |The Wheels Binding Point| $AN_2838 from movement(
  base_vel = {2.5},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA12:FSA(
            society[$AN_2852]<212,314>|State1| = [
              Stop]<100,100>
,
            society[$AN_2854]<476,171>|State2| = [
              CNP_BidOnTask]<100,100>
,
            society[$AN_2856]<748,314>|State3| = [
              Stop]<100,100>
,
            society[$AN_2858]<483,445>|State4| = [
              CNP_ExecuteWonTask]<100,100>
,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_2852,
            rules[$AN_2854]<476,171>|State2| = if [
              CNP_IsAuctionEnded]<0,0>|Trans1|
 goto $AN_2856,
            rules[$AN_2856]<748,314>|State3| = if [
              CNP_WonTask]<0,0>|Trans2|
 goto $AN_2858,
            rules[$AN_2856]<748,314>|State3| = if [
              CNP_LostTask]<0,0>|Trans3|
 goto $AN_2852,
            rules[$AN_2852]<212,314>|State1| = if [
              CNP_AuctionReady]<0,0>|Trans1|
 goto $AN_2854,
            rules[$AN_2858]<483,445>|State4| = if [
                %cnp_task = {CHECK_WON_CNP_TASK},
                %task_name = {""}
,
              CNP_TaskCompletionNotified]<335,374>|Trans1|
 goto $AN_2852)<292,156>|The State Machine|
,
        max_vel = {5.0},
        base_vel = {2.5},
        cautious_vel = {0.5},
        cautious_mode = {false})<222,15>|The Wheel Actuator|
);

instBP<100,100> $AN_2873 from vehicle(
  bound_to = sample-type-I-interceptRobot3:DEFAULT_ROBOT(
sample-type-I-interceptRobot3:[
          $AN_2838]
)<365,181>|Individual Robot|
);

instBP<222,15> |The Wheels Binding Point| $AN_2874 from movement(
  base_vel = {2.5},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA5:FSA(
            society[$AN_2852]<212,314>|State1| = [
              Stop]<100,100>
,
            society[$AN_2854]<476,171>|State2| = [
              CNP_BidOnTask]<100,100>
,
            society[$AN_2856]<748,314>|State3| = [
              Stop]<100,100>
,
            society[$AN_2858]<483,445>|State4| = [
              CNP_ExecuteWonTask]<100,100>
,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_2852,
            rules[$AN_2854]<476,171>|State2| = if [
              CNP_IsAuctionEnded]<0,0>|Trans1|
 goto $AN_2856,
            rules[$AN_2856]<748,314>|State3| = if [
              CNP_WonTask]<0,0>|Trans2|
 goto $AN_2858,
            rules[$AN_2856]<748,314>|State3| = if [
              CNP_LostTask]<0,0>|Trans3|
 goto $AN_2852,
            rules[$AN_2852]<212,314>|State1| = if [
              CNP_AuctionReady]<0,0>|Trans1|
 goto $AN_2854,
            rules[$AN_2858]<483,445>|State4| = if [
                %cnp_task = {CHECK_WON_CNP_TASK},
                %task_name = {""}
,
              CNP_TaskCompletionNotified]<335,374>|Trans1|
 goto $AN_2852)<292,156>|The State Machine|
,
        max_vel = {5.0},
        base_vel = {2.5},
        cautious_vel = {0.5},
        cautious_mode = {false})<222,15>|The Wheel Actuator|
);

instBP<100,100> $AN_2905 from vehicle(
  bound_to = sample-type-I-interceptRobot2:DEFAULT_ROBOT(
sample-type-I-interceptRobot2:[
          $AN_2874]
)<366,39>|Individual Robot|
);

instBP<222,15> |The Wheels Binding Point| $AN_2906 from movement(
  base_vel = {2.5},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA1:FSA(
            society[$AN_2960]<242,50>|State1| = [
              Stop]<10,10>
,
            society[$AN_2964]<240,222>|State2| = [
                %Objects = {Enemies}
,
              LookFor]<10,10>
,
            society[$AN_2968]<588,222>|State3| = [
                %Targets = {Enemy}
,
              CNP_SaveTargetLocation]<10,10>
,
            society[$AN_2972]<907,224>|State4| = [
                %Targets = {Enemy}
,
              CNP_SaveTargetVelocity]<10,10>
,
            society[$AN_2976]<906,446>|State5| = [
                %task_name = {"InterceptTask"},
                %task_id = {"0"},
                %task_constraints = {"ENVIRONMENT:0:SURFACE,MISSION_STEALTHINESS:0:NOT_STEALTHY,TARGET_LOCATION_X:2:*,TARGET_LOCATION_Y:2:*,TARGET_LOCATION_Z:2:*,TARGET_VELOCITY_X:2:*,TARGET_VELOCITY_Y:2:*,TARGET_VELOCITY_Z:2:*"}
,
              CNP_InjectTask]<10,10>
,
            society[$AN_2980]<597,448>|State6| = [
              Stop]<10,10>
,
            society[$AN_2984]<249,451>|State7| = [
                %alert_subject = {"Mission Accomplished"},
                %alert_message = {"The robot has completed all the tasks."},
                %sends_email = {NO_Email},
                %recipient = {""},
                %sends_image = {NO_Image}
,
              Alert]<10,10>
,
            society[Start]<50,50>|Start| = [
              Stop]<100,100>
,
            society[$AN_2996]<250,701>|State8| = [
              TerminateMission]<10,10>
,
            rules[$AN_2964]<240,222>|State2| = if [
                %Objects = {Enemies}
,
              Detect]<0,0>|Trans3|
 goto $AN_2968,
            rules[$AN_2968]<588,222>|State3| = if [
                %Delay = {2.0}
,
              Wait]<0,0>|Trans4|
 goto $AN_2972,
            rules[$AN_2972]<907,224>|State4| = if [
                %Delay = {2.0}
,
              Wait]<0,0>|Trans5|
 goto $AN_2976,
            rules[$AN_2976]<906,446>|State5| = if [
              Immediate]<0,0>|Trans6|
 goto $AN_2980,
            rules[$AN_2980]<597,448>|State6| = if [
                %cnp_task = {CHECK_SPECIFIC_CNP_TASK},
                %task_name = {"InterceptTask"}
,
              CNP_TaskCompletionNotified]<0,0>|Trans7|
 goto $AN_2984,
            rules[Start]<50,50>|Start| = if [
              Immediate]<0,0>|Trans1|
 goto $AN_2960,
            rules[$AN_2960]<242,50>|State1| = if [
                %Delay = {10.0}
,
              Wait]<0,0>|Trans2|
 goto $AN_2964,
            rules[$AN_2984]<249,451>|State7| = if [
              Alerted]<0,0>|Trans10|
 goto $AN_2996)<292,156>|The State Machine|
,
        max_vel = {5.0},
        base_vel = {2.5},
        cautious_vel = {0.5},
        cautious_mode = {false})<222,15>|The Wheel Actuator|
);

instBP<100,100> $AN_2957 from vehicle(
  bound_to = sample-type-I-interceptRobot1:DEFAULT_ROBOT(
sample-type-I-interceptRobot1:[
          $AN_2906]
)<49,38>|Individual Robot|
);

[
[
    $AN_2957,
    $AN_2905,
    $AN_2873]<10,10>|Group of Robots|
]<10,10>

