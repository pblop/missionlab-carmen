/*************************************************
*
* This CDL file sample_intercept.cdl was created with cfgedit
* version 6.0.01
*
**************************************************/

bindArch AuRA.naval;

instBP<222,15> |The Wheels Binding Point| $AN_2308 from movement(
  base_vel = {2.5},
  v<0,0> = ,
  bound_to = base:DRIVE_W_SPIN(
        v<12,15> = FSA1:FSA(
            society[Start]<50,50>|Start| = [
              Stop]<10,10>
,
            society[$AN_2323]<241,263>|State1| = [
              Stop]<10,10>
,
            society[$AN_2325]<663,262>|State2| = [
                %Objects = {Enemies},
                %intercept_gain = {1.0},
                %avoid_obstacle_gain = {0.5},
                %wander_gain = {0.0},
                %avoid_obstacle_sphere = {1.2},
                %avoid_obstacle_safety_margin = {0.3}
,
              Intercept]<10,10>
,
            society[$AN_2327]<665,492>|State3| = [
                %notify_message = {"Enemy stop."}
,
              NotifyRobots]<10,10>
,
            society[$AN_2329]<247,491>|State4| = [
              Stop]<10,10>
,
            rules[$AN_2323]<241,263>|State1| = if [
                %notify_message = {"Intercept."}
,
              Notified]<0,0>|Trans2|
 goto $AN_2325,
            rules[$AN_2325]<663,262>|State2| = if [
                %Objects = {Enemies},
                %Distance = {25.0}
,
              Near]<665,381>|Trans3|
 goto $AN_2327,
            rules[Start]<50,50>|Start| = if [
              Immediate]<10,10>|Trans1|
 goto $AN_2323,
            rules[$AN_2327]<665,492>|State3| = if [
              MessageSent]<10,10>|Trans5|
 goto $AN_2329)<292,156>|The State Machine|
,
        max_vel = {5.0},
        base_vel = {2.5},
        cautious_vel = {0.5},
        cautious_mode = {false})<222,15>|The Wheel Actuator|
);

instBP<0,0> $AN_2339 from vehicle(
  bound_to = sample_interceptRobot1:DEFAULT_ROBOT(
sample_interceptRobot1:[
          $AN_2308]
)<0,0>|Individual Robot|
);

[
[
    $AN_2339]<10,10>|Group of Robots|
]<10,10>

